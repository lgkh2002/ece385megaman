module metalman_rom (input [13:0] addr, output [3:0] data);




	parameter [0:9907][3:0] ROM = {
	
	
//	0: metal man standing
// 1: metal man pose 1
// 2: metal man pose 2
// 3: metal man run 1
// 4: metal man run 2
// 5: metal man run 3
// 6: metal man jump
// 7: metal throw 1
// 8: metal throw 2


//sawblade 1

4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd1,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,
4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd9,
4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,
4'd0,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd1,4'd0,4'd0,
4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,
4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,
4'd0,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd1,4'd0,4'd0,
4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,
4'd9,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,
4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd1,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,


//sawblade 2

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd9,4'd9,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd9,4'd9,
4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,
4'd9,4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd9,
4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,
4'd9,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd0,4'd9,
4'd9,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd0,4'd9,
4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,
4'd9,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,4'd9,
4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd1,4'd0,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd9,4'd9,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,






	
//metal man standing	
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd0,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,
	
	
	
	
//metal man pose 1

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd0,4'd3,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd3,4'd3,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd2,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd3,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd3,4'd3,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd0,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,


//metal man pose 2
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd3,4'd3,4'd0,4'd0,4'd2,4'd2,4'd0,4'd3,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd3,4'd2,4'd2,4'd2,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd0,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,	


//metal man run 1
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd3,4'd3,4'd3,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd3,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd2,4'd2,4'd0,4'd9,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,



//metal man run 2

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd2,4'd2,4'd0,4'd2,4'd2,4'd0,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,



//metal man run 3

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd3,4'd3,4'd2,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd3,4'd3,4'd3,4'd3,4'd3,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd3,4'd3,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
	
	

//metal man jump

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd9,4'd0,4'd2,4'd0,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd0,4'd2,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd9,4'd0,4'd0,4'd3,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd3,4'd3,4'd0,4'd3,4'd3,4'd3,4'd3,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd3,4'd3,4'd3,4'd3,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd3,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,	
	
	
	
//metal throw 1

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd1,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd2,4'd2,4'd2,4'd2,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd2,4'd0,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd3,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,	


//metal throw 2

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd1,4'd1,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd3,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd2,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd1,4'd2,4'd3,4'd3,4'd0,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd2,4'd3,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd1,4'd1,4'd1,4'd1,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd0,4'd2,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd0,4'd2,4'd3,4'd3,4'd0,4'd2,4'd2,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd0,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,
4'd9,4'd0,4'd2,4'd2,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd2,4'd2,4'd0,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd2,4'd2,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd2,4'd2,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd2,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9

	};

	assign data = ROM[addr];

endmodule 