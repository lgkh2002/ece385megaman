module megaman_rom ( input [13:0]	addr,
						output [2:0]	data
					 );

	parameter ADDR_WIDTH = 11;
   parameter DATA_WIDTH =  5;
	logic [ADDR_WIDTH-1:0] addr_reg;
	
	//2**ADDR_WIDTH-1
				
	// ROM definition				
	parameter [0:10277][2:0] ROM = {
	
	
	//0: standing - no gun
	//1: jumping - no gun 
	//2: run1 - no gun 
	//3: run2 - no gun 
	//4: run3 - no gun 
	//5: standing - with gun 
	//6: jumping - with gun
	//7: run1 - with gun
	//8: run2 - with gun
	//9: run3 - with gun
	//10: hurt
	
	
			//lemon
			3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,
			3'd5,3'd0,3'd6,3'd6,3'd6,3'd6,3'd0,3'd5,
			3'd0,3'd6,3'd6,3'd6,3'd4,3'd4,3'd6,3'd0,
			3'd0,3'd6,3'd6,3'd6,3'd6,3'd4,3'd6,3'd0,
			3'd5,3'd0,3'd6,3'd6,3'd6,3'd6,3'd0,3'd5,
			3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,
	
			
			
			//standing sprite
			
			//line 1
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			
			//line 2
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 3			
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 4						
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 5							
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 6
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			
			//line 7
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 8
			
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 9

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 10

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 11

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 12

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 13
			
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 14

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 13'd5,

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 16

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 17

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 18

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 19

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 20

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd2,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd2,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 21

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 22

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 23

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 24

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 23'd5,

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 26
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 27

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 28

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd0,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 29

			3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 30

			3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			
			//jumping sprite
			
			//line 3'd1,
			
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			
			//line 3'd2,
			
			3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 3'd3,
			
			3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,
			
			//line 3'd4,
			
			3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,
			
			//line 3'd5,
			
			3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,

			//line 6
			3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,

			//line 7 
			3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 8
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 9
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 10

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 11
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd0,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 12

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 13
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd3,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 14
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 15
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 16

			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 17
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 18
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 19
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,


			//line 20
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

			//line 21
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 22
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 23
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 24
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 25
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 26
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 27
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 28
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 29
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			
			//line 30
			3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
			

			//running sprite 1
			
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd0,3'd2,3'd2,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd5,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd0,3'd5,3'd0,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd0,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,


//running sprite 2

3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd2,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd2,3'd0,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd0,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd2,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,

	
//running sprite 3

3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd0,3'd1,3'd2,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd0,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5, 	
	
	
	
//standing with gun

3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd2,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd0,3'd2,3'd2,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd2,3'd0,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd2,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,	
	
	
	
	
//jump with gun

3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd2,3'd2,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd2,3'd0,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd0,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd3,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,	


//run 1 with gun

3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd0,3'd2,3'd2,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd2,3'd2,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd2,3'd0,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd5,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd0,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,


//run2 with gun

3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd2,3'd2,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd2,3'd0,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd2,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd2,3'd0,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd0,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd2,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,


//run3 with gun

3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd3,3'd4,3'd4,3'd0,3'd0,3'd3,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd2,3'd2,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd2,3'd0,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd1,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd0,3'd1,3'd2,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd0,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,


//hurt 
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd2,3'd2,3'd0,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd2,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd0,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd0,3'd2,3'd2,3'd0,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd0,3'd3,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,
3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd0,3'd0,3'd0,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5
	
        };

	assign data = ROM[addr];

endmodule  