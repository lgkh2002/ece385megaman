module enemy_rom(input [12:0] addr, output [3:0] data);


	parameter [0:4287][3:0] ROM = {
	
	//mole 1 (begins at 0) 8X24
	
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd5,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd3,4'd3,4'd0,4'd3,4'd3,4'd0,4'd8,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd0,4'd9,
4'd0,4'd7,4'd0,4'd7,4'd0,4'd7,4'd7,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd8,4'd0,
4'd0,4'd7,4'd0,4'd7,4'd0,4'd7,4'd7,4'd0,4'd5,4'd0,4'd5,4'd5,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd5,4'd0,4'd9,
4'd9,4'd0,4'd3,4'd3,4'd0,4'd3,4'd3,4'd0,4'd5,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd0,4'd8,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,

	//mole 2 (begins at 192) 8X24

4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd3,4'd3,4'd0,4'd3,4'd3,4'd0,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,
4'd0,4'd7,4'd0,4'd7,4'd0,4'd7,4'd7,4'd0,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd5,4'd8,4'd0,
4'd0,4'd7,4'd0,4'd7,4'd0,4'd7,4'd7,4'd0,4'd8,4'd5,4'd5,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd5,4'd0,4'd0,4'd9,
4'd9,4'd0,4'd3,4'd3,4'd0,4'd3,4'd3,4'd0,4'd8,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd8,4'd8,4'd0,4'd5,4'd8,4'd0,4'd5,4'd8,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,

	//pierobot 1 (begins at 384) 32X63
	
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd6,4'd6,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd6,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd6,4'd6,4'd6,4'd6,4'd4,4'd4,4'd0,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd6,4'd6,4'd4,4'd0,4'd9,4'd0,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd4,4'd4,4'd6,4'd0,4'd9,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd5,4'd5,4'd0,4'd0,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd5,4'd5,4'd0,4'd5,4'd5,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd5,4'd0,4'd5,4'd5,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd4,4'd4,4'd4,4'd0,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd5,4'd5,4'd4,4'd4,4'd0,4'd0,4'd4,4'd4,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd5,4'd0,4'd4,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd5,4'd5,4'd5,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd5,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd1,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd1,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd1,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd1,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd9,4'd9,
4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,
4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,
4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,
4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,
4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,
4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,
4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,
4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,
4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,
4'd9,4'd9,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd1,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd1,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd1,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd1,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,



// pierobot 2 (begins at 2368)

4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd3,4'd3,4'd3,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd6,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd6,4'd6,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd6,4'd6,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd6,4'd6,4'd6,4'd6,4'd6,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd1,4'd1,4'd0,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd5,4'd5,4'd0,4'd9,4'd0,4'd4,4'd0,4'd4,4'd0,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd5,4'd5,4'd0,4'd9,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd5,4'd0,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd5,4'd5,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd5,4'd5,4'd5,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd0,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd5,4'd5,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd1,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd1,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd1,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd1,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,
4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,
4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,
4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,
4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd1,4'd1,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd1,4'd1,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd1,4'd1,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd1,4'd1,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd9,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd9,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,
4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,

	
	};

	assign data = ROM[addr];

endmodule 